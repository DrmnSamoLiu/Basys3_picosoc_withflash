
module progmem
(
// Closk & reset
input  wire         clk,
input  wire         rstn,

// PicoRV32 bus interface
input  wire         valid,
output wire         ready,
input  wire [31:0]  addr,
output wire [31:0]  rdata
);

// ============================================================================

localparam  MEM_SIZE_BITS   = 11; // In 32-bit words
localparam  MEM_SIZE        = 1 << MEM_SIZE_BITS;
localparam  MEM_ADDR_MASK   = 32'h0010_0000;

// ============================================================================

wire [MEM_SIZE_BITS-1:0]    mem_addr;
reg  [31:0]                 mem_data;

always @(posedge clk)
    case (mem_addr)

    'h0000: mem_data <= 32'h00000093;
    'h0001: mem_data <= 32'h00000193;
    'h0002: mem_data <= 32'h00000213;
    'h0003: mem_data <= 32'h00000293;
    'h0004: mem_data <= 32'h00000313;
    'h0005: mem_data <= 32'h00000393;
    'h0006: mem_data <= 32'h00000413;
    'h0007: mem_data <= 32'h00000493;
    'h0008: mem_data <= 32'h00000513;
    'h0009: mem_data <= 32'h00000593;
    'h000A: mem_data <= 32'h00000613;
    'h000B: mem_data <= 32'h00000693;
    'h000C: mem_data <= 32'h00000713;
    'h000D: mem_data <= 32'h00000793;
    'h000E: mem_data <= 32'h00000813;
    'h000F: mem_data <= 32'h00000893;
    'h0010: mem_data <= 32'h00000913;
    'h0011: mem_data <= 32'h00000993;
    'h0012: mem_data <= 32'h00000A13;
    'h0013: mem_data <= 32'h00000A93;
    'h0014: mem_data <= 32'h00000B13;
    'h0015: mem_data <= 32'h00000B93;
    'h0016: mem_data <= 32'h00000C13;
    'h0017: mem_data <= 32'h00000C93;
    'h0018: mem_data <= 32'h00000D13;
    'h0019: mem_data <= 32'h00000D93;
    'h001A: mem_data <= 32'h00000E13;
    'h001B: mem_data <= 32'h00000E93;
    'h001C: mem_data <= 32'h00000F13;
    'h001D: mem_data <= 32'h00000F93;
    'h001E: mem_data <= 32'h03000537;
    'h001F: mem_data <= 32'h00100593;
    'h0020: mem_data <= 32'h00B52023;
    'h0021: mem_data <= 32'h00000513;
    'h0022: mem_data <= 32'h00A52023;
    'h0023: mem_data <= 32'h00450513;
    'h0024: mem_data <= 32'hFE254CE3;
    'h0025: mem_data <= 32'h03000537;
    'h0026: mem_data <= 32'h00300593;
    'h0027: mem_data <= 32'h00B52023;
    'h0028: mem_data <= 32'h00002517;
    'h0029: mem_data <= 32'hA6850513;
    'h002A: mem_data <= 32'h00000593;
    'h002B: mem_data <= 32'h00000613;
    'h002C: mem_data <= 32'h00C5DC63;
    'h002D: mem_data <= 32'h00052683;
    'h002E: mem_data <= 32'h00D5A023;
    'h002F: mem_data <= 32'h00450513;
    'h0030: mem_data <= 32'h00458593;
    'h0031: mem_data <= 32'hFEC5C8E3;
    'h0032: mem_data <= 32'h03000537;
    'h0033: mem_data <= 32'h00700593;
    'h0034: mem_data <= 32'h00B52023;
    'h0035: mem_data <= 32'h00000513;
    'h0036: mem_data <= 32'h00000593;
    'h0037: mem_data <= 32'h00B55863;
    'h0038: mem_data <= 32'h00052023;
    'h0039: mem_data <= 32'h00450513;
    'h003A: mem_data <= 32'hFEB54CE3;
    'h003B: mem_data <= 32'h03000537;
    'h003C: mem_data <= 32'h00F00593;
    'h003D: mem_data <= 32'h00B52023;
    'h003E: mem_data <= 32'h31C010EF;
    'h003F: mem_data <= 32'h0000006F;
    'h0040: mem_data <= 32'h020002B7;
    'h0041: mem_data <= 32'h12000313;
    'h0042: mem_data <= 32'h00629023;
    'h0043: mem_data <= 32'h000281A3;
    'h0044: mem_data <= 32'h02060863;
    'h0045: mem_data <= 32'h00800F13;
    'h0046: mem_data <= 32'h0FF67393;
    'h0047: mem_data <= 32'h0073DE93;
    'h0048: mem_data <= 32'h01D28023;
    'h0049: mem_data <= 32'h010EEE93;
    'h004A: mem_data <= 32'h01D28023;
    'h004B: mem_data <= 32'h00139393;
    'h004C: mem_data <= 32'h0FF3F393;
    'h004D: mem_data <= 32'hFFFF0F13;
    'h004E: mem_data <= 32'hFE0F12E3;
    'h004F: mem_data <= 32'h00628023;
    'h0050: mem_data <= 32'h04058663;
    'h0051: mem_data <= 32'h00800F13;
    'h0052: mem_data <= 32'h00054383;
    'h0053: mem_data <= 32'h0073DE93;
    'h0054: mem_data <= 32'h01D28023;
    'h0055: mem_data <= 32'h010EEE93;
    'h0056: mem_data <= 32'h01D28023;
    'h0057: mem_data <= 32'h0002CE83;
    'h0058: mem_data <= 32'h002EFE93;
    'h0059: mem_data <= 32'h001EDE93;
    'h005A: mem_data <= 32'h00139393;
    'h005B: mem_data <= 32'h01D3E3B3;
    'h005C: mem_data <= 32'h0FF3F393;
    'h005D: mem_data <= 32'hFFFF0F13;
    'h005E: mem_data <= 32'hFC0F1AE3;
    'h005F: mem_data <= 32'h00750023;
    'h0060: mem_data <= 32'h00150513;
    'h0061: mem_data <= 32'hFFF58593;
    'h0062: mem_data <= 32'hFB9FF06F;
    'h0063: mem_data <= 32'h08000313;
    'h0064: mem_data <= 32'h006281A3;
    'h0065: mem_data <= 32'h00008067;
    'h0066: mem_data <= 32'hFD010113;
    'h0067: mem_data <= 32'h02112623;
    'h0068: mem_data <= 32'h02812423;
    'h0069: mem_data <= 32'h02912223;
    'h006A: mem_data <= 32'h03010413;
    'h006B: mem_data <= 32'hFCA42E23;
    'h006C: mem_data <= 32'hFCB42C23;
    'h006D: mem_data <= 32'h00060693;
    'h006E: mem_data <= 32'hFCD40BA3;
    'h006F: mem_data <= 32'h00010693;
    'h0070: mem_data <= 32'h00068493;
    'h0071: mem_data <= 32'h001006B7;
    'h0072: mem_data <= 32'h19868613;
    'h0073: mem_data <= 32'h001006B7;
    'h0074: mem_data <= 32'h10068693;
    'h0075: mem_data <= 32'h40D606B3;
    'h0076: mem_data <= 32'h4026D693;
    'h0077: mem_data <= 32'hFFF68693;
    'h0078: mem_data <= 32'hFED42223;
    'h0079: mem_data <= 32'h001006B7;
    'h007A: mem_data <= 32'h19868613;
    'h007B: mem_data <= 32'h001006B7;
    'h007C: mem_data <= 32'h10068693;
    'h007D: mem_data <= 32'h40D606B3;
    'h007E: mem_data <= 32'h4026D693;
    'h007F: mem_data <= 32'h00068E13;
    'h0080: mem_data <= 32'h00000E93;
    'h0081: mem_data <= 32'h01BE5693;
    'h0082: mem_data <= 32'h005E9893;
    'h0083: mem_data <= 32'h0116E8B3;
    'h0084: mem_data <= 32'h005E1813;
    'h0085: mem_data <= 32'h001006B7;
    'h0086: mem_data <= 32'h19868613;
    'h0087: mem_data <= 32'h001006B7;
    'h0088: mem_data <= 32'h10068693;
    'h0089: mem_data <= 32'h40D606B3;
    'h008A: mem_data <= 32'h4026D693;
    'h008B: mem_data <= 32'h00068313;
    'h008C: mem_data <= 32'h00000393;
    'h008D: mem_data <= 32'h01B35693;
    'h008E: mem_data <= 32'h00539793;
    'h008F: mem_data <= 32'h00F6E7B3;
    'h0090: mem_data <= 32'h00531713;
    'h0091: mem_data <= 32'h001007B7;
    'h0092: mem_data <= 32'h19878713;
    'h0093: mem_data <= 32'h001007B7;
    'h0094: mem_data <= 32'h10078793;
    'h0095: mem_data <= 32'h40F707B3;
    'h0096: mem_data <= 32'h00378793;
    'h0097: mem_data <= 32'hFFC7F793;
    'h0098: mem_data <= 32'h00F78793;
    'h0099: mem_data <= 32'h0047D793;
    'h009A: mem_data <= 32'h00479793;
    'h009B: mem_data <= 32'h40F10133;
    'h009C: mem_data <= 32'h00010793;
    'h009D: mem_data <= 32'h00378793;
    'h009E: mem_data <= 32'h0027D793;
    'h009F: mem_data <= 32'h00279793;
    'h00A0: mem_data <= 32'hFEF42023;
    'h00A1: mem_data <= 32'h001007B7;
    'h00A2: mem_data <= 32'h10078793;
    'h00A3: mem_data <= 32'hFEF42423;
    'h00A4: mem_data <= 32'hFE042783;
    'h00A5: mem_data <= 32'hFEF42623;
    'h00A6: mem_data <= 32'h0240006F;
    'h00A7: mem_data <= 32'hFE842703;
    'h00A8: mem_data <= 32'h00470793;
    'h00A9: mem_data <= 32'hFEF42423;
    'h00AA: mem_data <= 32'hFEC42783;
    'h00AB: mem_data <= 32'h00478693;
    'h00AC: mem_data <= 32'hFED42623;
    'h00AD: mem_data <= 32'h00072703;
    'h00AE: mem_data <= 32'h00E7A023;
    'h00AF: mem_data <= 32'hFE842703;
    'h00B0: mem_data <= 32'h001007B7;
    'h00B1: mem_data <= 32'h19878793;
    'h00B2: mem_data <= 32'hFCF71AE3;
    'h00B3: mem_data <= 32'hFE042683;
    'h00B4: mem_data <= 32'hFD842783;
    'h00B5: mem_data <= 32'hFD744703;
    'h00B6: mem_data <= 32'h00070613;
    'h00B7: mem_data <= 32'h00078593;
    'h00B8: mem_data <= 32'hFDC42503;
    'h00B9: mem_data <= 32'h000680E7;
    'h00BA: mem_data <= 32'h00048113;
    'h00BB: mem_data <= 32'h00000013;
    'h00BC: mem_data <= 32'hFD040113;
    'h00BD: mem_data <= 32'h02C12083;
    'h00BE: mem_data <= 32'h02812403;
    'h00BF: mem_data <= 32'h02412483;
    'h00C0: mem_data <= 32'h03010113;
    'h00C1: mem_data <= 32'h00008067;
    'h00C2: mem_data <= 32'hFE010113;
    'h00C3: mem_data <= 32'h00112E23;
    'h00C4: mem_data <= 32'h00812C23;
    'h00C5: mem_data <= 32'h02010413;
    'h00C6: mem_data <= 32'h008007B7;
    'h00C7: mem_data <= 32'h00278793;
    'h00C8: mem_data <= 32'hFEF42623;
    'h00C9: mem_data <= 32'h06500793;
    'h00CA: mem_data <= 32'hFEF40023;
    'h00CB: mem_data <= 32'hFEC42783;
    'h00CC: mem_data <= 32'h0107D793;
    'h00CD: mem_data <= 32'h0FF7F793;
    'h00CE: mem_data <= 32'hFEF400A3;
    'h00CF: mem_data <= 32'hFEC42783;
    'h00D0: mem_data <= 32'h0087D793;
    'h00D1: mem_data <= 32'h0FF7F793;
    'h00D2: mem_data <= 32'hFEF40123;
    'h00D3: mem_data <= 32'hFEC42783;
    'h00D4: mem_data <= 32'h0FF7F793;
    'h00D5: mem_data <= 32'hFEF401A3;
    'h00D6: mem_data <= 32'hFE040223;
    'h00D7: mem_data <= 32'hFE0402A3;
    'h00D8: mem_data <= 32'hFE040793;
    'h00D9: mem_data <= 32'h00000613;
    'h00DA: mem_data <= 32'h00600593;
    'h00DB: mem_data <= 32'h00078513;
    'h00DC: mem_data <= 32'hE29FF0EF;
    'h00DD: mem_data <= 32'hFE544783;
    'h00DE: mem_data <= 32'hFEF405A3;
    'h00DF: mem_data <= 32'h07100793;
    'h00E0: mem_data <= 32'hFEF40023;
    'h00E1: mem_data <= 32'hFEC42783;
    'h00E2: mem_data <= 32'h0107D793;
    'h00E3: mem_data <= 32'h0FF7F793;
    'h00E4: mem_data <= 32'hFEF400A3;
    'h00E5: mem_data <= 32'hFEC42783;
    'h00E6: mem_data <= 32'h0087D793;
    'h00E7: mem_data <= 32'h0FF7F793;
    'h00E8: mem_data <= 32'hFEF40123;
    'h00E9: mem_data <= 32'hFEC42783;
    'h00EA: mem_data <= 32'h0FF7F793;
    'h00EB: mem_data <= 32'hFEF401A3;
    'h00EC: mem_data <= 32'hFEB44783;
    'h00ED: mem_data <= 32'h0027E793;
    'h00EE: mem_data <= 32'h0FF7F793;
    'h00EF: mem_data <= 32'hFEF40223;
    'h00F0: mem_data <= 32'hFE040793;
    'h00F1: mem_data <= 32'h00600613;
    'h00F2: mem_data <= 32'h00500593;
    'h00F3: mem_data <= 32'h00078513;
    'h00F4: mem_data <= 32'hDC9FF0EF;
    'h00F5: mem_data <= 32'h00000013;
    'h00F6: mem_data <= 32'h01C12083;
    'h00F7: mem_data <= 32'h01812403;
    'h00F8: mem_data <= 32'h02010113;
    'h00F9: mem_data <= 32'h00008067;
    'h00FA: mem_data <= 32'hFD010113;
    'h00FB: mem_data <= 32'h02112623;
    'h00FC: mem_data <= 32'h02812423;
    'h00FD: mem_data <= 32'h03010413;
    'h00FE: mem_data <= 32'h00050793;
    'h00FF: mem_data <= 32'hFCF40FA3;
    'h0100: mem_data <= 32'h020007B7;
    'h0101: mem_data <= 32'h0007A703;
    'h0102: mem_data <= 32'hFF8107B7;
    'h0103: mem_data <= 32'hFFF78793;
    'h0104: mem_data <= 32'h00F776B3;
    'h0105: mem_data <= 32'hFDF44783;
    'h0106: mem_data <= 32'h01079793;
    'h0107: mem_data <= 32'h00078713;
    'h0108: mem_data <= 32'h000F07B7;
    'h0109: mem_data <= 32'h00F77733;
    'h010A: mem_data <= 32'h020007B7;
    'h010B: mem_data <= 32'h00E6E733;
    'h010C: mem_data <= 32'h00E7A023;
    'h010D: mem_data <= 32'h008007B7;
    'h010E: mem_data <= 32'h00478793;
    'h010F: mem_data <= 32'hFEF42623;
    'h0110: mem_data <= 32'h07100793;
    'h0111: mem_data <= 32'hFEF40223;
    'h0112: mem_data <= 32'hFEC42783;
    'h0113: mem_data <= 32'h0107D793;
    'h0114: mem_data <= 32'h0FF7F793;
    'h0115: mem_data <= 32'hFEF402A3;
    'h0116: mem_data <= 32'hFEC42783;
    'h0117: mem_data <= 32'h0087D793;
    'h0118: mem_data <= 32'h0FF7F793;
    'h0119: mem_data <= 32'hFEF40323;
    'h011A: mem_data <= 32'hFEC42783;
    'h011B: mem_data <= 32'h0FF7F793;
    'h011C: mem_data <= 32'hFEF403A3;
    'h011D: mem_data <= 32'hFDF44783;
    'h011E: mem_data <= 32'h0707E793;
    'h011F: mem_data <= 32'h0FF7F793;
    'h0120: mem_data <= 32'hFEF40423;
    'h0121: mem_data <= 32'hFE440793;
    'h0122: mem_data <= 32'h00600613;
    'h0123: mem_data <= 32'h00500593;
    'h0124: mem_data <= 32'h00078513;
    'h0125: mem_data <= 32'hD05FF0EF;
    'h0126: mem_data <= 32'h00000013;
    'h0127: mem_data <= 32'h02C12083;
    'h0128: mem_data <= 32'h02812403;
    'h0129: mem_data <= 32'h03010113;
    'h012A: mem_data <= 32'h00008067;
    'h012B: mem_data <= 32'hFF010113;
    'h012C: mem_data <= 32'h00812623;
    'h012D: mem_data <= 32'h01010413;
    'h012E: mem_data <= 32'h020007B7;
    'h012F: mem_data <= 32'h0007A683;
    'h0130: mem_data <= 32'h020007B7;
    'h0131: mem_data <= 32'hFF900737;
    'h0132: mem_data <= 32'hFFF70713;
    'h0133: mem_data <= 32'h00E6F733;
    'h0134: mem_data <= 32'h00E7A023;
    'h0135: mem_data <= 32'h00000013;
    'h0136: mem_data <= 32'h00C12403;
    'h0137: mem_data <= 32'h01010113;
    'h0138: mem_data <= 32'h00008067;
    'h0139: mem_data <= 32'hFF010113;
    'h013A: mem_data <= 32'h00812623;
    'h013B: mem_data <= 32'h01010413;
    'h013C: mem_data <= 32'h020007B7;
    'h013D: mem_data <= 32'h0007A703;
    'h013E: mem_data <= 32'hFF9007B7;
    'h013F: mem_data <= 32'hFFF78793;
    'h0140: mem_data <= 32'h00F776B3;
    'h0141: mem_data <= 32'h020007B7;
    'h0142: mem_data <= 32'h00400737;
    'h0143: mem_data <= 32'h00E6E733;
    'h0144: mem_data <= 32'h00E7A023;
    'h0145: mem_data <= 32'h00000013;
    'h0146: mem_data <= 32'h00C12403;
    'h0147: mem_data <= 32'h01010113;
    'h0148: mem_data <= 32'h00008067;
    'h0149: mem_data <= 32'hFF010113;
    'h014A: mem_data <= 32'h00812623;
    'h014B: mem_data <= 32'h01010413;
    'h014C: mem_data <= 32'h020007B7;
    'h014D: mem_data <= 32'h0007A703;
    'h014E: mem_data <= 32'hFF9007B7;
    'h014F: mem_data <= 32'hFFF78793;
    'h0150: mem_data <= 32'h00F776B3;
    'h0151: mem_data <= 32'h020007B7;
    'h0152: mem_data <= 32'h00200737;
    'h0153: mem_data <= 32'h00E6E733;
    'h0154: mem_data <= 32'h00E7A023;
    'h0155: mem_data <= 32'h00000013;
    'h0156: mem_data <= 32'h00C12403;
    'h0157: mem_data <= 32'h01010113;
    'h0158: mem_data <= 32'h00008067;
    'h0159: mem_data <= 32'hFF010113;
    'h015A: mem_data <= 32'h00812623;
    'h015B: mem_data <= 32'h01010413;
    'h015C: mem_data <= 32'h020007B7;
    'h015D: mem_data <= 32'h0007A703;
    'h015E: mem_data <= 32'hFF9007B7;
    'h015F: mem_data <= 32'hFFF78793;
    'h0160: mem_data <= 32'h00F776B3;
    'h0161: mem_data <= 32'h020007B7;
    'h0162: mem_data <= 32'h00600737;
    'h0163: mem_data <= 32'h00E6E733;
    'h0164: mem_data <= 32'h00E7A023;
    'h0165: mem_data <= 32'h00000013;
    'h0166: mem_data <= 32'h00C12403;
    'h0167: mem_data <= 32'h01010113;
    'h0168: mem_data <= 32'h00008067;
    'h0169: mem_data <= 32'hFE010113;
    'h016A: mem_data <= 32'h00112E23;
    'h016B: mem_data <= 32'h00812C23;
    'h016C: mem_data <= 32'h02010413;
    'h016D: mem_data <= 32'h00050793;
    'h016E: mem_data <= 32'hFEF407A3;
    'h016F: mem_data <= 32'hFEF44703;
    'h0170: mem_data <= 32'h00A00793;
    'h0171: mem_data <= 32'h00F71663;
    'h0172: mem_data <= 32'h00D00513;
    'h0173: mem_data <= 32'hFD9FF0EF;
    'h0174: mem_data <= 32'h020007B7;
    'h0175: mem_data <= 32'h00878793;
    'h0176: mem_data <= 32'hFEF44703;
    'h0177: mem_data <= 32'h00E7A023;
    'h0178: mem_data <= 32'h00000013;
    'h0179: mem_data <= 32'h01C12083;
    'h017A: mem_data <= 32'h01812403;
    'h017B: mem_data <= 32'h02010113;
    'h017C: mem_data <= 32'h00008067;
    'h017D: mem_data <= 32'hFE010113;
    'h017E: mem_data <= 32'h00112E23;
    'h017F: mem_data <= 32'h00812C23;
    'h0180: mem_data <= 32'h02010413;
    'h0181: mem_data <= 32'hFEA42623;
    'h0182: mem_data <= 32'h01C0006F;
    'h0183: mem_data <= 32'hFEC42783;
    'h0184: mem_data <= 32'h00178713;
    'h0185: mem_data <= 32'hFEE42623;
    'h0186: mem_data <= 32'h0007C783;
    'h0187: mem_data <= 32'h00078513;
    'h0188: mem_data <= 32'hF85FF0EF;
    'h0189: mem_data <= 32'hFEC42783;
    'h018A: mem_data <= 32'h0007C783;
    'h018B: mem_data <= 32'hFE0790E3;
    'h018C: mem_data <= 32'h00000013;
    'h018D: mem_data <= 32'h00000013;
    'h018E: mem_data <= 32'h01C12083;
    'h018F: mem_data <= 32'h01812403;
    'h0190: mem_data <= 32'h02010113;
    'h0191: mem_data <= 32'h00008067;
    'h0192: mem_data <= 32'hFD010113;
    'h0193: mem_data <= 32'h02112623;
    'h0194: mem_data <= 32'h02812423;
    'h0195: mem_data <= 32'h03010413;
    'h0196: mem_data <= 32'hFCA42E23;
    'h0197: mem_data <= 32'hFCB42C23;
    'h0198: mem_data <= 32'h00700793;
    'h0199: mem_data <= 32'hFEF42623;
    'h019A: mem_data <= 32'h06C0006F;
    'h019B: mem_data <= 32'hFEC42783;
    'h019C: mem_data <= 32'h00279793;
    'h019D: mem_data <= 32'hFDC42703;
    'h019E: mem_data <= 32'h00F757B3;
    'h019F: mem_data <= 32'h00F7F793;
    'h01A0: mem_data <= 32'h00101737;
    'h01A1: mem_data <= 32'h77470713;
    'h01A2: mem_data <= 32'h00F707B3;
    'h01A3: mem_data <= 32'h0007C783;
    'h01A4: mem_data <= 32'hFEF405A3;
    'h01A5: mem_data <= 32'hFEB44703;
    'h01A6: mem_data <= 32'h03000793;
    'h01A7: mem_data <= 32'h00F71863;
    'h01A8: mem_data <= 32'hFEC42703;
    'h01A9: mem_data <= 32'hFD842783;
    'h01AA: mem_data <= 32'h00F75E63;
    'h01AB: mem_data <= 32'hFEB44783;
    'h01AC: mem_data <= 32'h00078513;
    'h01AD: mem_data <= 32'hEF1FF0EF;
    'h01AE: mem_data <= 32'hFEC42783;
    'h01AF: mem_data <= 32'hFCF42C23;
    'h01B0: mem_data <= 32'h0080006F;
    'h01B1: mem_data <= 32'h00000013;
    'h01B2: mem_data <= 32'hFEC42783;
    'h01B3: mem_data <= 32'hFFF78793;
    'h01B4: mem_data <= 32'hFEF42623;
    'h01B5: mem_data <= 32'hFEC42783;
    'h01B6: mem_data <= 32'hF807DAE3;
    'h01B7: mem_data <= 32'h00000013;
    'h01B8: mem_data <= 32'h00000013;
    'h01B9: mem_data <= 32'h02C12083;
    'h01BA: mem_data <= 32'h02812403;
    'h01BB: mem_data <= 32'h03010113;
    'h01BC: mem_data <= 32'h00008067;
    'h01BD: mem_data <= 32'hFE010113;
    'h01BE: mem_data <= 32'h00112E23;
    'h01BF: mem_data <= 32'h00812C23;
    'h01C0: mem_data <= 32'h02010413;
    'h01C1: mem_data <= 32'hFEA42623;
    'h01C2: mem_data <= 32'hFEC42703;
    'h01C3: mem_data <= 32'h06300793;
    'h01C4: mem_data <= 32'h00E7FA63;
    'h01C5: mem_data <= 32'h001017B7;
    'h01C6: mem_data <= 32'h78878513;
    'h01C7: mem_data <= 32'hED9FF0EF;
    'h01C8: mem_data <= 32'h28C0006F;
    'h01C9: mem_data <= 32'hFEC42703;
    'h01CA: mem_data <= 32'h05900793;
    'h01CB: mem_data <= 32'h00E7FE63;
    'h01CC: mem_data <= 32'h03900513;
    'h01CD: mem_data <= 32'hE71FF0EF;
    'h01CE: mem_data <= 32'hFEC42783;
    'h01CF: mem_data <= 32'hFA678793;
    'h01D0: mem_data <= 32'hFEF42623;
    'h01D1: mem_data <= 32'h1200006F;
    'h01D2: mem_data <= 32'hFEC42703;
    'h01D3: mem_data <= 32'h04F00793;
    'h01D4: mem_data <= 32'h00E7FE63;
    'h01D5: mem_data <= 32'h03800513;
    'h01D6: mem_data <= 32'hE4DFF0EF;
    'h01D7: mem_data <= 32'hFEC42783;
    'h01D8: mem_data <= 32'hFB078793;
    'h01D9: mem_data <= 32'hFEF42623;
    'h01DA: mem_data <= 32'h0FC0006F;
    'h01DB: mem_data <= 32'hFEC42703;
    'h01DC: mem_data <= 32'h04500793;
    'h01DD: mem_data <= 32'h00E7FE63;
    'h01DE: mem_data <= 32'h03700513;
    'h01DF: mem_data <= 32'hE29FF0EF;
    'h01E0: mem_data <= 32'hFEC42783;
    'h01E1: mem_data <= 32'hFBA78793;
    'h01E2: mem_data <= 32'hFEF42623;
    'h01E3: mem_data <= 32'h0D80006F;
    'h01E4: mem_data <= 32'hFEC42703;
    'h01E5: mem_data <= 32'h03B00793;
    'h01E6: mem_data <= 32'h00E7FE63;
    'h01E7: mem_data <= 32'h03600513;
    'h01E8: mem_data <= 32'hE05FF0EF;
    'h01E9: mem_data <= 32'hFEC42783;
    'h01EA: mem_data <= 32'hFC478793;
    'h01EB: mem_data <= 32'hFEF42623;
    'h01EC: mem_data <= 32'h0B40006F;
    'h01ED: mem_data <= 32'hFEC42703;
    'h01EE: mem_data <= 32'h03100793;
    'h01EF: mem_data <= 32'h00E7FE63;
    'h01F0: mem_data <= 32'h03500513;
    'h01F1: mem_data <= 32'hDE1FF0EF;
    'h01F2: mem_data <= 32'hFEC42783;
    'h01F3: mem_data <= 32'hFCE78793;
    'h01F4: mem_data <= 32'hFEF42623;
    'h01F5: mem_data <= 32'h0900006F;
    'h01F6: mem_data <= 32'hFEC42703;
    'h01F7: mem_data <= 32'h02700793;
    'h01F8: mem_data <= 32'h00E7FE63;
    'h01F9: mem_data <= 32'h03400513;
    'h01FA: mem_data <= 32'hDBDFF0EF;
    'h01FB: mem_data <= 32'hFEC42783;
    'h01FC: mem_data <= 32'hFD878793;
    'h01FD: mem_data <= 32'hFEF42623;
    'h01FE: mem_data <= 32'h06C0006F;
    'h01FF: mem_data <= 32'hFEC42703;
    'h0200: mem_data <= 32'h01D00793;
    'h0201: mem_data <= 32'h00E7FE63;
    'h0202: mem_data <= 32'h03300513;
    'h0203: mem_data <= 32'hD99FF0EF;
    'h0204: mem_data <= 32'hFEC42783;
    'h0205: mem_data <= 32'hFE278793;
    'h0206: mem_data <= 32'hFEF42623;
    'h0207: mem_data <= 32'h0480006F;
    'h0208: mem_data <= 32'hFEC42703;
    'h0209: mem_data <= 32'h01300793;
    'h020A: mem_data <= 32'h00E7FE63;
    'h020B: mem_data <= 32'h03200513;
    'h020C: mem_data <= 32'hD75FF0EF;
    'h020D: mem_data <= 32'hFEC42783;
    'h020E: mem_data <= 32'hFEC78793;
    'h020F: mem_data <= 32'hFEF42623;
    'h0210: mem_data <= 32'h0240006F;
    'h0211: mem_data <= 32'hFEC42703;
    'h0212: mem_data <= 32'h00900793;
    'h0213: mem_data <= 32'h00E7FC63;
    'h0214: mem_data <= 32'h03100513;
    'h0215: mem_data <= 32'hD51FF0EF;
    'h0216: mem_data <= 32'hFEC42783;
    'h0217: mem_data <= 32'hFF678793;
    'h0218: mem_data <= 32'hFEF42623;
    'h0219: mem_data <= 32'hFEC42703;
    'h021A: mem_data <= 32'h00800793;
    'h021B: mem_data <= 32'h00E7FE63;
    'h021C: mem_data <= 32'h03900513;
    'h021D: mem_data <= 32'hD31FF0EF;
    'h021E: mem_data <= 32'hFEC42783;
    'h021F: mem_data <= 32'hFF778793;
    'h0220: mem_data <= 32'hFEF42623;
    'h0221: mem_data <= 32'h1280006F;
    'h0222: mem_data <= 32'hFEC42703;
    'h0223: mem_data <= 32'h00700793;
    'h0224: mem_data <= 32'h00E7FE63;
    'h0225: mem_data <= 32'h03800513;
    'h0226: mem_data <= 32'hD0DFF0EF;
    'h0227: mem_data <= 32'hFEC42783;
    'h0228: mem_data <= 32'hFF878793;
    'h0229: mem_data <= 32'hFEF42623;
    'h022A: mem_data <= 32'h1040006F;
    'h022B: mem_data <= 32'hFEC42703;
    'h022C: mem_data <= 32'h00600793;
    'h022D: mem_data <= 32'h00E7FE63;
    'h022E: mem_data <= 32'h03700513;
    'h022F: mem_data <= 32'hCE9FF0EF;
    'h0230: mem_data <= 32'hFEC42783;
    'h0231: mem_data <= 32'hFF978793;
    'h0232: mem_data <= 32'hFEF42623;
    'h0233: mem_data <= 32'h0E00006F;
    'h0234: mem_data <= 32'hFEC42703;
    'h0235: mem_data <= 32'h00500793;
    'h0236: mem_data <= 32'h00E7FE63;
    'h0237: mem_data <= 32'h03600513;
    'h0238: mem_data <= 32'hCC5FF0EF;
    'h0239: mem_data <= 32'hFEC42783;
    'h023A: mem_data <= 32'hFFA78793;
    'h023B: mem_data <= 32'hFEF42623;
    'h023C: mem_data <= 32'h0BC0006F;
    'h023D: mem_data <= 32'hFEC42703;
    'h023E: mem_data <= 32'h00400793;
    'h023F: mem_data <= 32'h00E7FE63;
    'h0240: mem_data <= 32'h03500513;
    'h0241: mem_data <= 32'hCA1FF0EF;
    'h0242: mem_data <= 32'hFEC42783;
    'h0243: mem_data <= 32'hFFB78793;
    'h0244: mem_data <= 32'hFEF42623;
    'h0245: mem_data <= 32'h0980006F;
    'h0246: mem_data <= 32'hFEC42703;
    'h0247: mem_data <= 32'h00300793;
    'h0248: mem_data <= 32'h00E7FE63;
    'h0249: mem_data <= 32'h03400513;
    'h024A: mem_data <= 32'hC7DFF0EF;
    'h024B: mem_data <= 32'hFEC42783;
    'h024C: mem_data <= 32'hFFC78793;
    'h024D: mem_data <= 32'hFEF42623;
    'h024E: mem_data <= 32'h0740006F;
    'h024F: mem_data <= 32'hFEC42703;
    'h0250: mem_data <= 32'h00200793;
    'h0251: mem_data <= 32'h00E7FE63;
    'h0252: mem_data <= 32'h03300513;
    'h0253: mem_data <= 32'hC59FF0EF;
    'h0254: mem_data <= 32'hFEC42783;
    'h0255: mem_data <= 32'hFFD78793;
    'h0256: mem_data <= 32'hFEF42623;
    'h0257: mem_data <= 32'h0500006F;
    'h0258: mem_data <= 32'hFEC42703;
    'h0259: mem_data <= 32'h00100793;
    'h025A: mem_data <= 32'h00E7FE63;
    'h025B: mem_data <= 32'h03200513;
    'h025C: mem_data <= 32'hC35FF0EF;
    'h025D: mem_data <= 32'hFEC42783;
    'h025E: mem_data <= 32'hFFE78793;
    'h025F: mem_data <= 32'hFEF42623;
    'h0260: mem_data <= 32'h02C0006F;
    'h0261: mem_data <= 32'hFEC42783;
    'h0262: mem_data <= 32'h00078E63;
    'h0263: mem_data <= 32'h03100513;
    'h0264: mem_data <= 32'hC15FF0EF;
    'h0265: mem_data <= 32'hFEC42783;
    'h0266: mem_data <= 32'hFFF78793;
    'h0267: mem_data <= 32'hFEF42623;
    'h0268: mem_data <= 32'h00C0006F;
    'h0269: mem_data <= 32'h03000513;
    'h026A: mem_data <= 32'hBFDFF0EF;
    'h026B: mem_data <= 32'h01C12083;
    'h026C: mem_data <= 32'h01812403;
    'h026D: mem_data <= 32'h02010113;
    'h026E: mem_data <= 32'h00008067;
    'h026F: mem_data <= 32'hFD010113;
    'h0270: mem_data <= 32'h02112623;
    'h0271: mem_data <= 32'h02812423;
    'h0272: mem_data <= 32'h03010413;
    'h0273: mem_data <= 32'hFCA42E23;
    'h0274: mem_data <= 32'hFFF00793;
    'h0275: mem_data <= 32'hFEF42623;
    'h0276: mem_data <= 32'hC00027F3;
    'h0277: mem_data <= 32'hFEF42423;
    'h0278: mem_data <= 32'h030007B7;
    'h0279: mem_data <= 32'hFFF00713;
    'h027A: mem_data <= 32'h00E7A023;
    'h027B: mem_data <= 32'hFDC42783;
    'h027C: mem_data <= 32'h08078A63;
    'h027D: mem_data <= 32'hFDC42503;
    'h027E: mem_data <= 32'hBFDFF0EF;
    'h027F: mem_data <= 32'h0880006F;
    'h0280: mem_data <= 32'hC00027F3;
    'h0281: mem_data <= 32'hFEF42223;
    'h0282: mem_data <= 32'hFE442703;
    'h0283: mem_data <= 32'hFE842783;
    'h0284: mem_data <= 32'h40F707B3;
    'h0285: mem_data <= 32'hFEF42023;
    'h0286: mem_data <= 32'hFE042703;
    'h0287: mem_data <= 32'h00B727B7;
    'h0288: mem_data <= 32'hB0078793;
    'h0289: mem_data <= 32'h04E7F863;
    'h028A: mem_data <= 32'hFDC42783;
    'h028B: mem_data <= 32'h00078663;
    'h028C: mem_data <= 32'hFDC42503;
    'h028D: mem_data <= 32'hBC1FF0EF;
    'h028E: mem_data <= 32'hFE442783;
    'h028F: mem_data <= 32'hFEF42423;
    'h0290: mem_data <= 32'h030007B7;
    'h0291: mem_data <= 32'h0007A783;
    'h0292: mem_data <= 32'h00179713;
    'h0293: mem_data <= 32'h030007B7;
    'h0294: mem_data <= 32'h0007A783;
    'h0295: mem_data <= 32'h0017D793;
    'h0296: mem_data <= 32'h0017F793;
    'h0297: mem_data <= 32'h0017B793;
    'h0298: mem_data <= 32'h0FF7F793;
    'h0299: mem_data <= 32'h00078693;
    'h029A: mem_data <= 32'h030007B7;
    'h029B: mem_data <= 32'h00D76733;
    'h029C: mem_data <= 32'h00E7A023;
    'h029D: mem_data <= 32'h020007B7;
    'h029E: mem_data <= 32'h00878793;
    'h029F: mem_data <= 32'h0007A783;
    'h02A0: mem_data <= 32'hFEF42623;
    'h02A1: mem_data <= 32'hFEC42703;
    'h02A2: mem_data <= 32'hFFF00793;
    'h02A3: mem_data <= 32'hF6F70AE3;
    'h02A4: mem_data <= 32'h030007B7;
    'h02A5: mem_data <= 32'h0007A023;
    'h02A6: mem_data <= 32'hFEC42783;
    'h02A7: mem_data <= 32'h0FF7F793;
    'h02A8: mem_data <= 32'h00078513;
    'h02A9: mem_data <= 32'h02C12083;
    'h02AA: mem_data <= 32'h02812403;
    'h02AB: mem_data <= 32'h03010113;
    'h02AC: mem_data <= 32'h00008067;
    'h02AD: mem_data <= 32'hFF010113;
    'h02AE: mem_data <= 32'h00112623;
    'h02AF: mem_data <= 32'h00812423;
    'h02B0: mem_data <= 32'h01010413;
    'h02B1: mem_data <= 32'h00000513;
    'h02B2: mem_data <= 32'hEF5FF0EF;
    'h02B3: mem_data <= 32'h00050793;
    'h02B4: mem_data <= 32'h00078513;
    'h02B5: mem_data <= 32'h00C12083;
    'h02B6: mem_data <= 32'h00812403;
    'h02B7: mem_data <= 32'h01010113;
    'h02B8: mem_data <= 32'h00008067;
    'h02B9: mem_data <= 32'hFD010113;
    'h02BA: mem_data <= 32'h02112623;
    'h02BB: mem_data <= 32'h02812423;
    'h02BC: mem_data <= 32'h03010413;
    'h02BD: mem_data <= 32'h09F00793;
    'h02BE: mem_data <= 32'hFCF42C23;
    'h02BF: mem_data <= 32'hFC042E23;
    'h02C0: mem_data <= 32'hFE042023;
    'h02C1: mem_data <= 32'hFE042223;
    'h02C2: mem_data <= 32'hFE040423;
    'h02C3: mem_data <= 32'hFD840793;
    'h02C4: mem_data <= 32'h00000613;
    'h02C5: mem_data <= 32'h01100593;
    'h02C6: mem_data <= 32'h00078513;
    'h02C7: mem_data <= 32'hE7CFF0EF;
    'h02C8: mem_data <= 32'h00100793;
    'h02C9: mem_data <= 32'hFEF42623;
    'h02CA: mem_data <= 32'h0340006F;
    'h02CB: mem_data <= 32'h02000513;
    'h02CC: mem_data <= 32'hA75FF0EF;
    'h02CD: mem_data <= 32'hFEC42783;
    'h02CE: mem_data <= 32'hFF040713;
    'h02CF: mem_data <= 32'h00F707B3;
    'h02D0: mem_data <= 32'hFE87C783;
    'h02D1: mem_data <= 32'h00200593;
    'h02D2: mem_data <= 32'h00078513;
    'h02D3: mem_data <= 32'hAFDFF0EF;
    'h02D4: mem_data <= 32'hFEC42783;
    'h02D5: mem_data <= 32'h00178793;
    'h02D6: mem_data <= 32'hFEF42623;
    'h02D7: mem_data <= 32'hFEC42703;
    'h02D8: mem_data <= 32'h01000793;
    'h02D9: mem_data <= 32'hFCE7D4E3;
    'h02DA: mem_data <= 32'h00A00513;
    'h02DB: mem_data <= 32'hA39FF0EF;
    'h02DC: mem_data <= 32'h00000013;
    'h02DD: mem_data <= 32'h02C12083;
    'h02DE: mem_data <= 32'h02812403;
    'h02DF: mem_data <= 32'h03010113;
    'h02E0: mem_data <= 32'h00008067;
    'h02E1: mem_data <= 32'hFD010113;
    'h02E2: mem_data <= 32'h02112623;
    'h02E3: mem_data <= 32'h02812423;
    'h02E4: mem_data <= 32'h03010413;
    'h02E5: mem_data <= 32'hFCA42E23;
    'h02E6: mem_data <= 32'hFCB42C23;
    'h02E7: mem_data <= 32'h00800513;
    'h02E8: mem_data <= 32'h849FF0EF;
    'h02E9: mem_data <= 32'h06500793;
    'h02EA: mem_data <= 32'hFEF40423;
    'h02EB: mem_data <= 32'hFDC42783;
    'h02EC: mem_data <= 32'h0107D793;
    'h02ED: mem_data <= 32'h0FF7F793;
    'h02EE: mem_data <= 32'hFEF404A3;
    'h02EF: mem_data <= 32'hFDC42783;
    'h02F0: mem_data <= 32'h0087D793;
    'h02F1: mem_data <= 32'h0FF7F793;
    'h02F2: mem_data <= 32'hFEF40523;
    'h02F3: mem_data <= 32'hFDC42783;
    'h02F4: mem_data <= 32'h0FF7F793;
    'h02F5: mem_data <= 32'hFEF405A3;
    'h02F6: mem_data <= 32'hFE040623;
    'h02F7: mem_data <= 32'hFE0406A3;
    'h02F8: mem_data <= 32'hFE840793;
    'h02F9: mem_data <= 32'h00000613;
    'h02FA: mem_data <= 32'h00600593;
    'h02FB: mem_data <= 32'h00078513;
    'h02FC: mem_data <= 32'hDA8FF0EF;
    'h02FD: mem_data <= 32'h001017B7;
    'h02FE: mem_data <= 32'h79078513;
    'h02FF: mem_data <= 32'h9F9FF0EF;
    'h0300: mem_data <= 32'h00600593;
    'h0301: mem_data <= 32'hFDC42503;
    'h0302: mem_data <= 32'hA41FF0EF;
    'h0303: mem_data <= 32'h001017B7;
    'h0304: mem_data <= 32'h79478513;
    'h0305: mem_data <= 32'h9E1FF0EF;
    'h0306: mem_data <= 32'hFD842503;
    'h0307: mem_data <= 32'h9D9FF0EF;
    'h0308: mem_data <= 32'h001017B7;
    'h0309: mem_data <= 32'h79878513;
    'h030A: mem_data <= 32'h9CDFF0EF;
    'h030B: mem_data <= 32'hFED44783;
    'h030C: mem_data <= 32'h00200593;
    'h030D: mem_data <= 32'h00078513;
    'h030E: mem_data <= 32'hA11FF0EF;
    'h030F: mem_data <= 32'h001017B7;
    'h0310: mem_data <= 32'h79C78513;
    'h0311: mem_data <= 32'h9B1FF0EF;
    'h0312: mem_data <= 32'hFED44783;
    'h0313: mem_data <= 32'h00078513;
    'h0314: mem_data <= 32'h02C12083;
    'h0315: mem_data <= 32'h02812403;
    'h0316: mem_data <= 32'h03010113;
    'h0317: mem_data <= 32'h00008067;
    'h0318: mem_data <= 32'hFE010113;
    'h0319: mem_data <= 32'h00112E23;
    'h031A: mem_data <= 32'h00812C23;
    'h031B: mem_data <= 32'h02010413;
    'h031C: mem_data <= 32'h001017B7;
    'h031D: mem_data <= 32'h79C78513;
    'h031E: mem_data <= 32'h97DFF0EF;
    'h031F: mem_data <= 32'h001017B7;
    'h0320: mem_data <= 32'h7A078593;
    'h0321: mem_data <= 32'h00800537;
    'h0322: mem_data <= 32'hEFDFF0EF;
    'h0323: mem_data <= 32'h00050793;
    'h0324: mem_data <= 32'hFEF407A3;
    'h0325: mem_data <= 32'h001017B7;
    'h0326: mem_data <= 32'h7A878593;
    'h0327: mem_data <= 32'h008007B7;
    'h0328: mem_data <= 32'h00178513;
    'h0329: mem_data <= 32'hEE1FF0EF;
    'h032A: mem_data <= 32'h00050793;
    'h032B: mem_data <= 32'hFEF40723;
    'h032C: mem_data <= 32'h001017B7;
    'h032D: mem_data <= 32'h7B078593;
    'h032E: mem_data <= 32'h008007B7;
    'h032F: mem_data <= 32'h00278513;
    'h0330: mem_data <= 32'hEC5FF0EF;
    'h0331: mem_data <= 32'h00050793;
    'h0332: mem_data <= 32'hFEF406A3;
    'h0333: mem_data <= 32'h001017B7;
    'h0334: mem_data <= 32'h7B878593;
    'h0335: mem_data <= 32'h008007B7;
    'h0336: mem_data <= 32'h00378513;
    'h0337: mem_data <= 32'hEA9FF0EF;
    'h0338: mem_data <= 32'h00050793;
    'h0339: mem_data <= 32'hFEF40623;
    'h033A: mem_data <= 32'h001017B7;
    'h033B: mem_data <= 32'h7C078593;
    'h033C: mem_data <= 32'h008007B7;
    'h033D: mem_data <= 32'h00478513;
    'h033E: mem_data <= 32'hE8DFF0EF;
    'h033F: mem_data <= 32'h00050793;
    'h0340: mem_data <= 32'hFEF405A3;
    'h0341: mem_data <= 32'h001017B7;
    'h0342: mem_data <= 32'h7C878593;
    'h0343: mem_data <= 32'h008007B7;
    'h0344: mem_data <= 32'h00578513;
    'h0345: mem_data <= 32'hE71FF0EF;
    'h0346: mem_data <= 32'h00050793;
    'h0347: mem_data <= 32'hFEF40523;
    'h0348: mem_data <= 32'h00000013;
    'h0349: mem_data <= 32'h01C12083;
    'h034A: mem_data <= 32'h01812403;
    'h034B: mem_data <= 32'h02010113;
    'h034C: mem_data <= 32'h00008067;
    'h034D: mem_data <= 32'hEB010113;
    'h034E: mem_data <= 32'h14112623;
    'h034F: mem_data <= 32'h14812423;
    'h0350: mem_data <= 32'h15010413;
    'h0351: mem_data <= 32'h00050793;
    'h0352: mem_data <= 32'hEAB42C23;
    'h0353: mem_data <= 32'hEAF40FA3;
    'h0354: mem_data <= 32'hEC040793;
    'h0355: mem_data <= 32'hFCF42A23;
    'h0356: mem_data <= 32'h12B9B7B7;
    'h0357: mem_data <= 32'h0A178793;
    'h0358: mem_data <= 32'hFEF42623;
    'h0359: mem_data <= 32'hC00027F3;
    'h035A: mem_data <= 32'hFCF42823;
    'h035B: mem_data <= 32'hC02027F3;
    'h035C: mem_data <= 32'hFCF42623;
    'h035D: mem_data <= 32'hFE042423;
    'h035E: mem_data <= 32'h1200006F;
    'h035F: mem_data <= 32'hFE042223;
    'h0360: mem_data <= 32'h0640006F;
    'h0361: mem_data <= 32'hFEC42783;
    'h0362: mem_data <= 32'h00D79793;
    'h0363: mem_data <= 32'hFEC42703;
    'h0364: mem_data <= 32'h00F747B3;
    'h0365: mem_data <= 32'hFEF42623;
    'h0366: mem_data <= 32'hFEC42783;
    'h0367: mem_data <= 32'h0117D793;
    'h0368: mem_data <= 32'hFEC42703;
    'h0369: mem_data <= 32'h00F747B3;
    'h036A: mem_data <= 32'hFEF42623;
    'h036B: mem_data <= 32'hFEC42783;
    'h036C: mem_data <= 32'h00579793;
    'h036D: mem_data <= 32'hFEC42703;
    'h036E: mem_data <= 32'h00F747B3;
    'h036F: mem_data <= 32'hFEF42623;
    'h0370: mem_data <= 32'hFEC42783;
    'h0371: mem_data <= 32'h0FF7F713;
    'h0372: mem_data <= 32'hFE442783;
    'h0373: mem_data <= 32'hFF040693;
    'h0374: mem_data <= 32'h00F687B3;
    'h0375: mem_data <= 32'hECE78823;
    'h0376: mem_data <= 32'hFE442783;
    'h0377: mem_data <= 32'h00178793;
    'h0378: mem_data <= 32'hFEF42223;
    'h0379: mem_data <= 32'hFE442703;
    'h037A: mem_data <= 32'h0FF00793;
    'h037B: mem_data <= 32'hF8E7DCE3;
    'h037C: mem_data <= 32'hFE042023;
    'h037D: mem_data <= 32'hFC042E23;
    'h037E: mem_data <= 32'h0440006F;
    'h037F: mem_data <= 32'hFE042783;
    'h0380: mem_data <= 32'hFF040713;
    'h0381: mem_data <= 32'h00F707B3;
    'h0382: mem_data <= 32'hED07C783;
    'h0383: mem_data <= 32'h02078263;
    'h0384: mem_data <= 32'hFDC42783;
    'h0385: mem_data <= 32'h00178713;
    'h0386: mem_data <= 32'hFCE42E23;
    'h0387: mem_data <= 32'hFE042703;
    'h0388: mem_data <= 32'h0FF77713;
    'h0389: mem_data <= 32'hFF040693;
    'h038A: mem_data <= 32'h00F687B3;
    'h038B: mem_data <= 32'hECE78823;
    'h038C: mem_data <= 32'hFE042783;
    'h038D: mem_data <= 32'h00178793;
    'h038E: mem_data <= 32'hFEF42023;
    'h038F: mem_data <= 32'hFE042703;
    'h0390: mem_data <= 32'h0FF00793;
    'h0391: mem_data <= 32'hFAE7DCE3;
    'h0392: mem_data <= 32'hFC042C23;
    'h0393: mem_data <= 32'hFC042023;
    'h0394: mem_data <= 32'h0300006F;
    'h0395: mem_data <= 32'hFD842783;
    'h0396: mem_data <= 32'h00279793;
    'h0397: mem_data <= 32'hFD442703;
    'h0398: mem_data <= 32'h00F707B3;
    'h0399: mem_data <= 32'h0007A783;
    'h039A: mem_data <= 32'hFEC42703;
    'h039B: mem_data <= 32'h00F747B3;
    'h039C: mem_data <= 32'hFEF42623;
    'h039D: mem_data <= 32'hFD842783;
    'h039E: mem_data <= 32'h00178793;
    'h039F: mem_data <= 32'hFCF42C23;
    'h03A0: mem_data <= 32'hFD842703;
    'h03A1: mem_data <= 32'h03F00793;
    'h03A2: mem_data <= 32'hFCE7D6E3;
    'h03A3: mem_data <= 32'hFE842783;
    'h03A4: mem_data <= 32'h00178793;
    'h03A5: mem_data <= 32'hFEF42423;
    'h03A6: mem_data <= 32'hFE842703;
    'h03A7: mem_data <= 32'h01300793;
    'h03A8: mem_data <= 32'hECE7DEE3;
    'h03A9: mem_data <= 32'hC00027F3;
    'h03AA: mem_data <= 32'hFCF42423;
    'h03AB: mem_data <= 32'hC02027F3;
    'h03AC: mem_data <= 32'hFCF42223;
    'h03AD: mem_data <= 32'hEBF44783;
    'h03AE: mem_data <= 32'h06078E63;
    'h03AF: mem_data <= 32'h001017B7;
    'h03B0: mem_data <= 32'h7D078513;
    'h03B1: mem_data <= 32'hF30FF0EF;
    'h03B2: mem_data <= 32'hFC842703;
    'h03B3: mem_data <= 32'hFD042783;
    'h03B4: mem_data <= 32'h40F707B3;
    'h03B5: mem_data <= 32'h00800593;
    'h03B6: mem_data <= 32'h00078513;
    'h03B7: mem_data <= 32'hF6CFF0EF;
    'h03B8: mem_data <= 32'h00A00513;
    'h03B9: mem_data <= 32'hEC0FF0EF;
    'h03BA: mem_data <= 32'h001017B7;
    'h03BB: mem_data <= 32'h7DC78513;
    'h03BC: mem_data <= 32'hF04FF0EF;
    'h03BD: mem_data <= 32'hFC442703;
    'h03BE: mem_data <= 32'hFCC42783;
    'h03BF: mem_data <= 32'h40F707B3;
    'h03C0: mem_data <= 32'h00800593;
    'h03C1: mem_data <= 32'h00078513;
    'h03C2: mem_data <= 32'hF40FF0EF;
    'h03C3: mem_data <= 32'h00A00513;
    'h03C4: mem_data <= 32'hE94FF0EF;
    'h03C5: mem_data <= 32'h001017B7;
    'h03C6: mem_data <= 32'h7E878513;
    'h03C7: mem_data <= 32'hED8FF0EF;
    'h03C8: mem_data <= 32'h00800593;
    'h03C9: mem_data <= 32'hFEC42503;
    'h03CA: mem_data <= 32'hF20FF0EF;
    'h03CB: mem_data <= 32'h00A00513;
    'h03CC: mem_data <= 32'hE74FF0EF;
    'h03CD: mem_data <= 32'hEB842783;
    'h03CE: mem_data <= 32'h00078C63;
    'h03CF: mem_data <= 32'hFC442703;
    'h03D0: mem_data <= 32'hFCC42783;
    'h03D1: mem_data <= 32'h40F70733;
    'h03D2: mem_data <= 32'hEB842783;
    'h03D3: mem_data <= 32'h00E7A023;
    'h03D4: mem_data <= 32'hFC842703;
    'h03D5: mem_data <= 32'hFD042783;
    'h03D6: mem_data <= 32'h40F707B3;
    'h03D7: mem_data <= 32'h00078513;
    'h03D8: mem_data <= 32'h14C12083;
    'h03D9: mem_data <= 32'h14812403;
    'h03DA: mem_data <= 32'h15010113;
    'h03DB: mem_data <= 32'h00008067;
    'h03DC: mem_data <= 32'hFD010113;
    'h03DD: mem_data <= 32'h02112623;
    'h03DE: mem_data <= 32'h02812423;
    'h03DF: mem_data <= 32'h03010413;
    'h03E0: mem_data <= 32'hFC042A23;
    'h03E1: mem_data <= 32'h001017B7;
    'h03E2: mem_data <= 32'h7F478513;
    'h03E3: mem_data <= 32'hE68FF0EF;
    'h03E4: mem_data <= 32'h020007B7;
    'h03E5: mem_data <= 32'h0007A683;
    'h03E6: mem_data <= 32'h020007B7;
    'h03E7: mem_data <= 32'hFF900737;
    'h03E8: mem_data <= 32'hFFF70713;
    'h03E9: mem_data <= 32'h00E6F733;
    'h03EA: mem_data <= 32'h00E7A023;
    'h03EB: mem_data <= 32'h001027B7;
    'h03EC: mem_data <= 32'h80478513;
    'h03ED: mem_data <= 32'hE40FF0EF;
    'h03EE: mem_data <= 32'hFD440793;
    'h03EF: mem_data <= 32'h00078593;
    'h03F0: mem_data <= 32'h00000513;
    'h03F1: mem_data <= 32'hD71FF0EF;
    'h03F2: mem_data <= 32'h00050793;
    'h03F3: mem_data <= 32'h00800593;
    'h03F4: mem_data <= 32'h00078513;
    'h03F5: mem_data <= 32'hE74FF0EF;
    'h03F6: mem_data <= 32'h00A00513;
    'h03F7: mem_data <= 32'hDC8FF0EF;
    'h03F8: mem_data <= 32'h00800793;
    'h03F9: mem_data <= 32'hFEF42623;
    'h03FA: mem_data <= 32'h09C0006F;
    'h03FB: mem_data <= 32'h001027B7;
    'h03FC: mem_data <= 32'h80878513;
    'h03FD: mem_data <= 32'hE00FF0EF;
    'h03FE: mem_data <= 32'hFEC42783;
    'h03FF: mem_data <= 32'h00078513;
    'h0400: mem_data <= 32'hEF4FF0EF;
    'h0401: mem_data <= 32'h001027B7;
    'h0402: mem_data <= 32'h81078513;
    'h0403: mem_data <= 32'hDE8FF0EF;
    'h0404: mem_data <= 32'hFEC42783;
    'h0405: mem_data <= 32'h0FF7F793;
    'h0406: mem_data <= 32'h00078513;
    'h0407: mem_data <= 32'hBCCFF0EF;
    'h0408: mem_data <= 32'h020007B7;
    'h0409: mem_data <= 32'h0007A703;
    'h040A: mem_data <= 32'hFF9007B7;
    'h040B: mem_data <= 32'hFFF78793;
    'h040C: mem_data <= 32'h00F776B3;
    'h040D: mem_data <= 32'h020007B7;
    'h040E: mem_data <= 32'h00400737;
    'h040F: mem_data <= 32'h00E6E733;
    'h0410: mem_data <= 32'h00E7A023;
    'h0411: mem_data <= 32'h001027B7;
    'h0412: mem_data <= 32'h80478513;
    'h0413: mem_data <= 32'hDA8FF0EF;
    'h0414: mem_data <= 32'hFD440793;
    'h0415: mem_data <= 32'h00078593;
    'h0416: mem_data <= 32'h00000513;
    'h0417: mem_data <= 32'hCD9FF0EF;
    'h0418: mem_data <= 32'h00050793;
    'h0419: mem_data <= 32'h00800593;
    'h041A: mem_data <= 32'h00078513;
    'h041B: mem_data <= 32'hDDCFF0EF;
    'h041C: mem_data <= 32'h00A00513;
    'h041D: mem_data <= 32'hD30FF0EF;
    'h041E: mem_data <= 32'hFEC42783;
    'h041F: mem_data <= 32'hFFF78793;
    'h0420: mem_data <= 32'hFEF42623;
    'h0421: mem_data <= 32'hFEC42783;
    'h0422: mem_data <= 32'hF6F042E3;
    'h0423: mem_data <= 32'h00800793;
    'h0424: mem_data <= 32'hFEF42423;
    'h0425: mem_data <= 32'h09C0006F;
    'h0426: mem_data <= 32'h001027B7;
    'h0427: mem_data <= 32'h81C78513;
    'h0428: mem_data <= 32'hD54FF0EF;
    'h0429: mem_data <= 32'hFE842783;
    'h042A: mem_data <= 32'h00078513;
    'h042B: mem_data <= 32'hE48FF0EF;
    'h042C: mem_data <= 32'h001027B7;
    'h042D: mem_data <= 32'h82878513;
    'h042E: mem_data <= 32'hD3CFF0EF;
    'h042F: mem_data <= 32'hFE842783;
    'h0430: mem_data <= 32'h0FF7F793;
    'h0431: mem_data <= 32'h00078513;
    'h0432: mem_data <= 32'hB20FF0EF;
    'h0433: mem_data <= 32'h020007B7;
    'h0434: mem_data <= 32'h0007A703;
    'h0435: mem_data <= 32'hFF9007B7;
    'h0436: mem_data <= 32'hFFF78793;
    'h0437: mem_data <= 32'h00F776B3;
    'h0438: mem_data <= 32'h020007B7;
    'h0439: mem_data <= 32'h00500737;
    'h043A: mem_data <= 32'h00E6E733;
    'h043B: mem_data <= 32'h00E7A023;
    'h043C: mem_data <= 32'h001027B7;
    'h043D: mem_data <= 32'h80478513;
    'h043E: mem_data <= 32'hCFCFF0EF;
    'h043F: mem_data <= 32'hFD440793;
    'h0440: mem_data <= 32'h00078593;
    'h0441: mem_data <= 32'h00000513;
    'h0442: mem_data <= 32'hC2DFF0EF;
    'h0443: mem_data <= 32'h00050793;
    'h0444: mem_data <= 32'h00800593;
    'h0445: mem_data <= 32'h00078513;
    'h0446: mem_data <= 32'hD30FF0EF;
    'h0447: mem_data <= 32'h00A00513;
    'h0448: mem_data <= 32'hC84FF0EF;
    'h0449: mem_data <= 32'hFE842783;
    'h044A: mem_data <= 32'hFFF78793;
    'h044B: mem_data <= 32'hFEF42423;
    'h044C: mem_data <= 32'hFE842783;
    'h044D: mem_data <= 32'hF6F042E3;
    'h044E: mem_data <= 32'h00800793;
    'h044F: mem_data <= 32'hFEF42223;
    'h0450: mem_data <= 32'h09C0006F;
    'h0451: mem_data <= 32'h001027B7;
    'h0452: mem_data <= 32'h83078513;
    'h0453: mem_data <= 32'hCA8FF0EF;
    'h0454: mem_data <= 32'hFE442783;
    'h0455: mem_data <= 32'h00078513;
    'h0456: mem_data <= 32'hD9CFF0EF;
    'h0457: mem_data <= 32'h001027B7;
    'h0458: mem_data <= 32'h81078513;
    'h0459: mem_data <= 32'hC90FF0EF;
    'h045A: mem_data <= 32'hFE442783;
    'h045B: mem_data <= 32'h0FF7F793;
    'h045C: mem_data <= 32'h00078513;
    'h045D: mem_data <= 32'hA74FF0EF;
    'h045E: mem_data <= 32'h020007B7;
    'h045F: mem_data <= 32'h0007A703;
    'h0460: mem_data <= 32'hFF9007B7;
    'h0461: mem_data <= 32'hFFF78793;
    'h0462: mem_data <= 32'h00F776B3;
    'h0463: mem_data <= 32'h020007B7;
    'h0464: mem_data <= 32'h00200737;
    'h0465: mem_data <= 32'h00E6E733;
    'h0466: mem_data <= 32'h00E7A023;
    'h0467: mem_data <= 32'h001027B7;
    'h0468: mem_data <= 32'h80478513;
    'h0469: mem_data <= 32'hC50FF0EF;
    'h046A: mem_data <= 32'hFD440793;
    'h046B: mem_data <= 32'h00078593;
    'h046C: mem_data <= 32'h00000513;
    'h046D: mem_data <= 32'hB81FF0EF;
    'h046E: mem_data <= 32'h00050793;
    'h046F: mem_data <= 32'h00800593;
    'h0470: mem_data <= 32'h00078513;
    'h0471: mem_data <= 32'hC84FF0EF;
    'h0472: mem_data <= 32'h00A00513;
    'h0473: mem_data <= 32'hBD8FF0EF;
    'h0474: mem_data <= 32'hFE442783;
    'h0475: mem_data <= 32'hFFF78793;
    'h0476: mem_data <= 32'hFEF42223;
    'h0477: mem_data <= 32'hFE442783;
    'h0478: mem_data <= 32'hF6F042E3;
    'h0479: mem_data <= 32'h00800793;
    'h047A: mem_data <= 32'hFEF42023;
    'h047B: mem_data <= 32'h09C0006F;
    'h047C: mem_data <= 32'h001027B7;
    'h047D: mem_data <= 32'h83878513;
    'h047E: mem_data <= 32'hBFCFF0EF;
    'h047F: mem_data <= 32'hFE042783;
    'h0480: mem_data <= 32'h00078513;
    'h0481: mem_data <= 32'hCF0FF0EF;
    'h0482: mem_data <= 32'h001027B7;
    'h0483: mem_data <= 32'h82878513;
    'h0484: mem_data <= 32'hBE4FF0EF;
    'h0485: mem_data <= 32'hFE042783;
    'h0486: mem_data <= 32'h0FF7F793;
    'h0487: mem_data <= 32'h00078513;
    'h0488: mem_data <= 32'h9C8FF0EF;
    'h0489: mem_data <= 32'h020007B7;
    'h048A: mem_data <= 32'h0007A703;
    'h048B: mem_data <= 32'hFF9007B7;
    'h048C: mem_data <= 32'hFFF78793;
    'h048D: mem_data <= 32'h00F776B3;
    'h048E: mem_data <= 32'h020007B7;
    'h048F: mem_data <= 32'h00300737;
    'h0490: mem_data <= 32'h00E6E733;
    'h0491: mem_data <= 32'h00E7A023;
    'h0492: mem_data <= 32'h001027B7;
    'h0493: mem_data <= 32'h80478513;
    'h0494: mem_data <= 32'hBA4FF0EF;
    'h0495: mem_data <= 32'hFD440793;
    'h0496: mem_data <= 32'h00078593;
    'h0497: mem_data <= 32'h00000513;
    'h0498: mem_data <= 32'hAD5FF0EF;
    'h0499: mem_data <= 32'h00050793;
    'h049A: mem_data <= 32'h00800593;
    'h049B: mem_data <= 32'h00078513;
    'h049C: mem_data <= 32'hBD8FF0EF;
    'h049D: mem_data <= 32'h00A00513;
    'h049E: mem_data <= 32'hB2CFF0EF;
    'h049F: mem_data <= 32'hFE042783;
    'h04A0: mem_data <= 32'hFFF78793;
    'h04A1: mem_data <= 32'hFEF42023;
    'h04A2: mem_data <= 32'hFE042783;
    'h04A3: mem_data <= 32'hF6F042E3;
    'h04A4: mem_data <= 32'h00800793;
    'h04A5: mem_data <= 32'hFCF42E23;
    'h04A6: mem_data <= 32'h09C0006F;
    'h04A7: mem_data <= 32'h001027B7;
    'h04A8: mem_data <= 32'h84478513;
    'h04A9: mem_data <= 32'hB50FF0EF;
    'h04AA: mem_data <= 32'hFDC42783;
    'h04AB: mem_data <= 32'h00078513;
    'h04AC: mem_data <= 32'hC44FF0EF;
    'h04AD: mem_data <= 32'h001027B7;
    'h04AE: mem_data <= 32'h82878513;
    'h04AF: mem_data <= 32'hB38FF0EF;
    'h04B0: mem_data <= 32'hFDC42783;
    'h04B1: mem_data <= 32'h0FF7F793;
    'h04B2: mem_data <= 32'h00078513;
    'h04B3: mem_data <= 32'h91CFF0EF;
    'h04B4: mem_data <= 32'h020007B7;
    'h04B5: mem_data <= 32'h0007A703;
    'h04B6: mem_data <= 32'hFF9007B7;
    'h04B7: mem_data <= 32'hFFF78793;
    'h04B8: mem_data <= 32'h00F776B3;
    'h04B9: mem_data <= 32'h020007B7;
    'h04BA: mem_data <= 32'h00600737;
    'h04BB: mem_data <= 32'h00E6E733;
    'h04BC: mem_data <= 32'h00E7A023;
    'h04BD: mem_data <= 32'h001027B7;
    'h04BE: mem_data <= 32'h80478513;
    'h04BF: mem_data <= 32'hAF8FF0EF;
    'h04C0: mem_data <= 32'hFD440793;
    'h04C1: mem_data <= 32'h00078593;
    'h04C2: mem_data <= 32'h00000513;
    'h04C3: mem_data <= 32'hA29FF0EF;
    'h04C4: mem_data <= 32'h00050793;
    'h04C5: mem_data <= 32'h00800593;
    'h04C6: mem_data <= 32'h00078513;
    'h04C7: mem_data <= 32'hB2CFF0EF;
    'h04C8: mem_data <= 32'h00A00513;
    'h04C9: mem_data <= 32'hA80FF0EF;
    'h04CA: mem_data <= 32'hFDC42783;
    'h04CB: mem_data <= 32'hFFF78793;
    'h04CC: mem_data <= 32'hFCF42E23;
    'h04CD: mem_data <= 32'hFDC42783;
    'h04CE: mem_data <= 32'hF6F042E3;
    'h04CF: mem_data <= 32'h00800793;
    'h04D0: mem_data <= 32'hFCF42C23;
    'h04D1: mem_data <= 32'h0900006F;
    'h04D2: mem_data <= 32'h001027B7;
    'h04D3: mem_data <= 32'h85078513;
    'h04D4: mem_data <= 32'hAA4FF0EF;
    'h04D5: mem_data <= 32'hFD842783;
    'h04D6: mem_data <= 32'h00078513;
    'h04D7: mem_data <= 32'hB98FF0EF;
    'h04D8: mem_data <= 32'h001017B7;
    'h04D9: mem_data <= 32'h79478513;
    'h04DA: mem_data <= 32'hA8CFF0EF;
    'h04DB: mem_data <= 32'hFD842783;
    'h04DC: mem_data <= 32'h0FF7F793;
    'h04DD: mem_data <= 32'h00078513;
    'h04DE: mem_data <= 32'h870FF0EF;
    'h04DF: mem_data <= 32'h020007B7;
    'h04E0: mem_data <= 32'h0007A683;
    'h04E1: mem_data <= 32'h020007B7;
    'h04E2: mem_data <= 32'h00700737;
    'h04E3: mem_data <= 32'h00E6E733;
    'h04E4: mem_data <= 32'h00E7A023;
    'h04E5: mem_data <= 32'h001027B7;
    'h04E6: mem_data <= 32'h80478513;
    'h04E7: mem_data <= 32'hA58FF0EF;
    'h04E8: mem_data <= 32'hFD440793;
    'h04E9: mem_data <= 32'h00078593;
    'h04EA: mem_data <= 32'h00000513;
    'h04EB: mem_data <= 32'h989FF0EF;
    'h04EC: mem_data <= 32'h00050793;
    'h04ED: mem_data <= 32'h00800593;
    'h04EE: mem_data <= 32'h00078513;
    'h04EF: mem_data <= 32'hA8CFF0EF;
    'h04F0: mem_data <= 32'h00A00513;
    'h04F1: mem_data <= 32'h9E0FF0EF;
    'h04F2: mem_data <= 32'hFD842783;
    'h04F3: mem_data <= 32'hFFF78793;
    'h04F4: mem_data <= 32'hFCF42C23;
    'h04F5: mem_data <= 32'hFD842783;
    'h04F6: mem_data <= 32'hF6F048E3;
    'h04F7: mem_data <= 32'h001027B7;
    'h04F8: mem_data <= 32'h86078513;
    'h04F9: mem_data <= 32'hA10FF0EF;
    'h04FA: mem_data <= 32'hFD442783;
    'h04FB: mem_data <= 32'h00800593;
    'h04FC: mem_data <= 32'h00078513;
    'h04FD: mem_data <= 32'hA54FF0EF;
    'h04FE: mem_data <= 32'h00A00513;
    'h04FF: mem_data <= 32'h9A8FF0EF;
    'h0500: mem_data <= 32'h00000013;
    'h0501: mem_data <= 32'h02C12083;
    'h0502: mem_data <= 32'h02812403;
    'h0503: mem_data <= 32'h03010113;
    'h0504: mem_data <= 32'h00008067;
    'h0505: mem_data <= 32'hFE010113;
    'h0506: mem_data <= 32'h00112E23;
    'h0507: mem_data <= 32'h00812C23;
    'h0508: mem_data <= 32'h02010413;
    'h0509: mem_data <= 32'h030007B7;
    'h050A: mem_data <= 32'h01F00713;
    'h050B: mem_data <= 32'h00E7A023;
    'h050C: mem_data <= 32'h020007B7;
    'h050D: mem_data <= 32'h00478793;
    'h050E: mem_data <= 32'h36400713;
    'h050F: mem_data <= 32'h00E7A023;
    'h0510: mem_data <= 32'h001027B7;
    'h0511: mem_data <= 32'h87478513;
    'h0512: mem_data <= 32'h9ACFF0EF;
    'h0513: mem_data <= 32'h030007B7;
    'h0514: mem_data <= 32'h03F00713;
    'h0515: mem_data <= 32'h00E7A023;
    'h0516: mem_data <= 32'hEB1FE0EF;
    'h0517: mem_data <= 32'h030007B7;
    'h0518: mem_data <= 32'h07F00713;
    'h0519: mem_data <= 32'h00E7A023;
    'h051A: mem_data <= 32'h00000013;
    'h051B: mem_data <= 32'h001027B7;
    'h051C: mem_data <= 32'h88078513;
    'h051D: mem_data <= 32'hD48FF0EF;
    'h051E: mem_data <= 32'h00050793;
    'h051F: mem_data <= 32'h00078713;
    'h0520: mem_data <= 32'h00D00793;
    'h0521: mem_data <= 32'hFEF714E3;
    'h0522: mem_data <= 32'h001017B7;
    'h0523: mem_data <= 32'h79C78513;
    'h0524: mem_data <= 32'h964FF0EF;
    'h0525: mem_data <= 32'h001027B7;
    'h0526: mem_data <= 32'h89C78513;
    'h0527: mem_data <= 32'h958FF0EF;
    'h0528: mem_data <= 32'h001027B7;
    'h0529: mem_data <= 32'h8C478513;
    'h052A: mem_data <= 32'h94CFF0EF;
    'h052B: mem_data <= 32'h001027B7;
    'h052C: mem_data <= 32'h8EC78513;
    'h052D: mem_data <= 32'h940FF0EF;
    'h052E: mem_data <= 32'h001027B7;
    'h052F: mem_data <= 32'h91078513;
    'h0530: mem_data <= 32'h934FF0EF;
    'h0531: mem_data <= 32'h001027B7;
    'h0532: mem_data <= 32'h93878513;
    'h0533: mem_data <= 32'h928FF0EF;
    'h0534: mem_data <= 32'h001017B7;
    'h0535: mem_data <= 32'h79C78513;
    'h0536: mem_data <= 32'h91CFF0EF;
    'h0537: mem_data <= 32'h001017B7;
    'h0538: mem_data <= 32'h79C78513;
    'h0539: mem_data <= 32'h910FF0EF;
    'h053A: mem_data <= 32'h001027B7;
    'h053B: mem_data <= 32'h96078513;
    'h053C: mem_data <= 32'h904FF0EF;
    'h053D: mem_data <= 32'h001027B7;
    'h053E: mem_data <= 32'h96C78513;
    'h053F: mem_data <= 32'h8F8FF0EF;
    'h0540: mem_data <= 32'h020007B7;
    'h0541: mem_data <= 32'h0007A783;
    'h0542: mem_data <= 32'h0107D793;
    'h0543: mem_data <= 32'h00F7F793;
    'h0544: mem_data <= 32'h00078513;
    'h0545: mem_data <= 32'h9E0FF0EF;
    'h0546: mem_data <= 32'h001017B7;
    'h0547: mem_data <= 32'h79C78513;
    'h0548: mem_data <= 32'h8D4FF0EF;
    'h0549: mem_data <= 32'h001027B7;
    'h054A: mem_data <= 32'h97878513;
    'h054B: mem_data <= 32'h8C8FF0EF;
    'h054C: mem_data <= 32'h020007B7;
    'h054D: mem_data <= 32'h0007A703;
    'h054E: mem_data <= 32'h004007B7;
    'h054F: mem_data <= 32'h00F777B3;
    'h0550: mem_data <= 32'h00078A63;
    'h0551: mem_data <= 32'h001027B7;
    'h0552: mem_data <= 32'h98078513;
    'h0553: mem_data <= 32'h8A8FF0EF;
    'h0554: mem_data <= 32'h0100006F;
    'h0555: mem_data <= 32'h001027B7;
    'h0556: mem_data <= 32'h98478513;
    'h0557: mem_data <= 32'h898FF0EF;
    'h0558: mem_data <= 32'h001027B7;
    'h0559: mem_data <= 32'h98C78513;
    'h055A: mem_data <= 32'h88CFF0EF;
    'h055B: mem_data <= 32'h020007B7;
    'h055C: mem_data <= 32'h0007A703;
    'h055D: mem_data <= 32'h002007B7;
    'h055E: mem_data <= 32'h00F777B3;
    'h055F: mem_data <= 32'h00078A63;
    'h0560: mem_data <= 32'h001027B7;
    'h0561: mem_data <= 32'h98078513;
    'h0562: mem_data <= 32'h86CFF0EF;
    'h0563: mem_data <= 32'h0100006F;
    'h0564: mem_data <= 32'h001027B7;
    'h0565: mem_data <= 32'h98478513;
    'h0566: mem_data <= 32'h85CFF0EF;
    'h0567: mem_data <= 32'h001027B7;
    'h0568: mem_data <= 32'h99478513;
    'h0569: mem_data <= 32'h850FF0EF;
    'h056A: mem_data <= 32'h020007B7;
    'h056B: mem_data <= 32'h0007A703;
    'h056C: mem_data <= 32'h001007B7;
    'h056D: mem_data <= 32'h00F777B3;
    'h056E: mem_data <= 32'h00078A63;
    'h056F: mem_data <= 32'h001027B7;
    'h0570: mem_data <= 32'h98078513;
    'h0571: mem_data <= 32'h830FF0EF;
    'h0572: mem_data <= 32'h0100006F;
    'h0573: mem_data <= 32'h001027B7;
    'h0574: mem_data <= 32'h98478513;
    'h0575: mem_data <= 32'h820FF0EF;
    'h0576: mem_data <= 32'h001017B7;
    'h0577: mem_data <= 32'h79C78513;
    'h0578: mem_data <= 32'h814FF0EF;
    'h0579: mem_data <= 32'h001027B7;
    'h057A: mem_data <= 32'h99C78513;
    'h057B: mem_data <= 32'h808FF0EF;
    'h057C: mem_data <= 32'h001017B7;
    'h057D: mem_data <= 32'h79C78513;
    'h057E: mem_data <= 32'hFFDFE0EF;
    'h057F: mem_data <= 32'h001027B7;
    'h0580: mem_data <= 32'h9B078513;
    'h0581: mem_data <= 32'hFF1FE0EF;
    'h0582: mem_data <= 32'h001027B7;
    'h0583: mem_data <= 32'h9CC78513;
    'h0584: mem_data <= 32'hFE5FE0EF;
    'h0585: mem_data <= 32'h001027B7;
    'h0586: mem_data <= 32'h9EC78513;
    'h0587: mem_data <= 32'hFD9FE0EF;
    'h0588: mem_data <= 32'h001027B7;
    'h0589: mem_data <= 32'hA0C78513;
    'h058A: mem_data <= 32'hFCDFE0EF;
    'h058B: mem_data <= 32'h001027B7;
    'h058C: mem_data <= 32'hA2C78513;
    'h058D: mem_data <= 32'hFC1FE0EF;
    'h058E: mem_data <= 32'h001027B7;
    'h058F: mem_data <= 32'hA4C78513;
    'h0590: mem_data <= 32'hFB5FE0EF;
    'h0591: mem_data <= 32'h001027B7;
    'h0592: mem_data <= 32'hA6C78513;
    'h0593: mem_data <= 32'hFA9FE0EF;
    'h0594: mem_data <= 32'h001027B7;
    'h0595: mem_data <= 32'hA9078513;
    'h0596: mem_data <= 32'hF9DFE0EF;
    'h0597: mem_data <= 32'h001027B7;
    'h0598: mem_data <= 32'hAB478513;
    'h0599: mem_data <= 32'hF91FE0EF;
    'h059A: mem_data <= 32'h001017B7;
    'h059B: mem_data <= 32'h79C78513;
    'h059C: mem_data <= 32'hF85FE0EF;
    'h059D: mem_data <= 32'h00A00793;
    'h059E: mem_data <= 32'hFEF42623;
    'h059F: mem_data <= 32'h0EC0006F;
    'h05A0: mem_data <= 32'h001027B7;
    'h05A1: mem_data <= 32'hAD478513;
    'h05A2: mem_data <= 32'hF6DFE0EF;
    'h05A3: mem_data <= 32'hC28FF0EF;
    'h05A4: mem_data <= 32'h00050793;
    'h05A5: mem_data <= 32'hFEF405A3;
    'h05A6: mem_data <= 32'hFEB44703;
    'h05A7: mem_data <= 32'h02000793;
    'h05A8: mem_data <= 32'h00E7FE63;
    'h05A9: mem_data <= 32'hFEB44703;
    'h05AA: mem_data <= 32'h07E00793;
    'h05AB: mem_data <= 32'h00E7E863;
    'h05AC: mem_data <= 32'hFEB44783;
    'h05AD: mem_data <= 32'h00078513;
    'h05AE: mem_data <= 32'hEEDFE0EF;
    'h05AF: mem_data <= 32'h001017B7;
    'h05B0: mem_data <= 32'h79C78513;
    'h05B1: mem_data <= 32'hF31FE0EF;
    'h05B2: mem_data <= 32'hFEB44783;
    'h05B3: mem_data <= 32'hFD078793;
    'h05B4: mem_data <= 32'h00900713;
    'h05B5: mem_data <= 32'h08F76063;
    'h05B6: mem_data <= 32'h00279713;
    'h05B7: mem_data <= 32'h001027B7;
    'h05B8: mem_data <= 32'hAE078793;
    'h05B9: mem_data <= 32'h00F707B3;
    'h05BA: mem_data <= 32'h0007A783;
    'h05BB: mem_data <= 32'h00078067;
    'h05BC: mem_data <= 32'hBF4FF0EF;
    'h05BD: mem_data <= 32'h0700006F;
    'h05BE: mem_data <= 32'hD68FF0EF;
    'h05BF: mem_data <= 32'h0680006F;
    'h05C0: mem_data <= 32'hDADFE0EF;
    'h05C1: mem_data <= 32'h0600006F;
    'h05C2: mem_data <= 32'hDDDFE0EF;
    'h05C3: mem_data <= 32'h0580006F;
    'h05C4: mem_data <= 32'hE15FE0EF;
    'h05C5: mem_data <= 32'h0500006F;
    'h05C6: mem_data <= 32'hE4DFE0EF;
    'h05C7: mem_data <= 32'h0480006F;
    'h05C8: mem_data <= 32'h020007B7;
    'h05C9: mem_data <= 32'h0007A683;
    'h05CA: mem_data <= 32'h020007B7;
    'h05CB: mem_data <= 32'h00100737;
    'h05CC: mem_data <= 32'h00E6C733;
    'h05CD: mem_data <= 32'h00E7A023;
    'h05CE: mem_data <= 32'h02C0006F;
    'h05CF: mem_data <= 32'h00000593;
    'h05D0: mem_data <= 32'h00100513;
    'h05D1: mem_data <= 32'hDF0FF0EF;
    'h05D2: mem_data <= 32'h01C0006F;
    'h05D3: mem_data <= 32'h825FF0EF;
    'h05D4: mem_data <= 32'h0140006F;
    'h05D5: mem_data <= 32'hFEC42783;
    'h05D6: mem_data <= 32'hFFF78793;
    'h05D7: mem_data <= 32'hFEF42623;
    'h05D8: mem_data <= 32'h0080006F;
    'h05D9: mem_data <= 32'h00C0006F;
    'h05DA: mem_data <= 32'hFEC42783;
    'h05DB: mem_data <= 32'hF0F04AE3;
    'h05DC: mem_data <= 32'hD61FF06F;
    'h05DD: mem_data <= 32'h33323130;
    'h05DE: mem_data <= 32'h37363534;
    'h05DF: mem_data <= 32'h62613938;
    'h05E0: mem_data <= 32'h66656463;
    'h05E1: mem_data <= 32'h00000000;
    'h05E2: mem_data <= 32'h30313D3E;
    'h05E3: mem_data <= 32'h00000030;
    'h05E4: mem_data <= 32'h00007830;
    'h05E5: mem_data <= 32'h00000020;
    'h05E6: mem_data <= 32'h00783020;
    'h05E7: mem_data <= 32'h0000000A;
    'h05E8: mem_data <= 32'h56315253;
    'h05E9: mem_data <= 32'h00000000;
    'h05EA: mem_data <= 32'h56325253;
    'h05EB: mem_data <= 32'h00000000;
    'h05EC: mem_data <= 32'h56315243;
    'h05ED: mem_data <= 32'h00000000;
    'h05EE: mem_data <= 32'h56325243;
    'h05EF: mem_data <= 32'h00000000;
    'h05F0: mem_data <= 32'h56335243;
    'h05F1: mem_data <= 32'h00000000;
    'h05F2: mem_data <= 32'h504C4456;
    'h05F3: mem_data <= 32'h00000000;
    'h05F4: mem_data <= 32'h6C637943;
    'h05F5: mem_data <= 32'h203A7365;
    'h05F6: mem_data <= 32'h00007830;
    'h05F7: mem_data <= 32'h74736E49;
    'h05F8: mem_data <= 32'h203A736E;
    'h05F9: mem_data <= 32'h00007830;
    'h05FA: mem_data <= 32'h736B6843;
    'h05FB: mem_data <= 32'h203A6D75;
    'h05FC: mem_data <= 32'h00007830;
    'h05FD: mem_data <= 32'h61666564;
    'h05FE: mem_data <= 32'h20746C75;
    'h05FF: mem_data <= 32'h20202020;
    'h0600: mem_data <= 32'h00202020;
    'h0601: mem_data <= 32'h0000203A;
    'h0602: mem_data <= 32'h69707364;
    'h0603: mem_data <= 32'h0000002D;
    'h0604: mem_data <= 32'h20202020;
    'h0605: mem_data <= 32'h20202020;
    'h0606: mem_data <= 32'h00000020;
    'h0607: mem_data <= 32'h69707364;
    'h0608: mem_data <= 32'h6D72632D;
    'h0609: mem_data <= 32'h0000002D;
    'h060A: mem_data <= 32'h20202020;
    'h060B: mem_data <= 32'h00000020;
    'h060C: mem_data <= 32'h69707371;
    'h060D: mem_data <= 32'h0000002D;
    'h060E: mem_data <= 32'h69707371;
    'h060F: mem_data <= 32'h6D72632D;
    'h0610: mem_data <= 32'h0000002D;
    'h0611: mem_data <= 32'h69707371;
    'h0612: mem_data <= 32'h7264642D;
    'h0613: mem_data <= 32'h0000002D;
    'h0614: mem_data <= 32'h69707371;
    'h0615: mem_data <= 32'h7264642D;
    'h0616: mem_data <= 32'h6D72632D;
    'h0617: mem_data <= 32'h0000002D;
    'h0618: mem_data <= 32'h74736E69;
    'h0619: mem_data <= 32'h2020736E;
    'h061A: mem_data <= 32'h20202020;
    'h061B: mem_data <= 32'h3A202020;
    'h061C: mem_data <= 32'h00000020;
    'h061D: mem_data <= 32'h746F6F42;
    'h061E: mem_data <= 32'h2E676E69;
    'h061F: mem_data <= 32'h00000A2E;
    'h0620: mem_data <= 32'h73657250;
    'h0621: mem_data <= 32'h4E452073;
    'h0622: mem_data <= 32'h20524554;
    'h0623: mem_data <= 32'h63206F74;
    'h0624: mem_data <= 32'h69746E6F;
    'h0625: mem_data <= 32'h2E65756E;
    'h0626: mem_data <= 32'h00000A2E;
    'h0627: mem_data <= 32'h5F5F2020;
    'h0628: mem_data <= 32'h20205F5F;
    'h0629: mem_data <= 32'h2020205F;
    'h062A: mem_data <= 32'h20202020;
    'h062B: mem_data <= 32'h5F202020;
    'h062C: mem_data <= 32'h205F5F5F;
    'h062D: mem_data <= 32'h20202020;
    'h062E: mem_data <= 32'h20202020;
    'h062F: mem_data <= 32'h5F5F5F5F;
    'h0630: mem_data <= 32'h0000000A;
    'h0631: mem_data <= 32'h20207C20;
    'h0632: mem_data <= 32'h285C205F;
    'h0633: mem_data <= 32'h5F20295F;
    'h0634: mem_data <= 32'h5F205F5F;
    'h0635: mem_data <= 32'h202F5F5F;
    'h0636: mem_data <= 32'h7C5F5F5F;
    'h0637: mem_data <= 32'h5F5F2020;
    'h0638: mem_data <= 32'h2F20205F;
    'h0639: mem_data <= 32'h5F5F5F20;
    'h063A: mem_data <= 32'h00000A7C;
    'h063B: mem_data <= 32'h7C207C20;
    'h063C: mem_data <= 32'h7C20295F;
    'h063D: mem_data <= 32'h202F7C20;
    'h063E: mem_data <= 32'h202F5F5F;
    'h063F: mem_data <= 32'h5F5C205F;
    'h0640: mem_data <= 32'h5C205F5F;
    'h0641: mem_data <= 32'h5F202F20;
    'h0642: mem_data <= 32'h207C5C20;
    'h0643: mem_data <= 32'h00000A7C;
    'h0644: mem_data <= 32'h20207C20;
    'h0645: mem_data <= 32'h7C2F5F5F;
    'h0646: mem_data <= 32'h28207C20;
    'h0647: mem_data <= 32'h28207C5F;
    'h0648: mem_data <= 32'h7C20295F;
    'h0649: mem_data <= 32'h20295F5F;
    'h064A: mem_data <= 32'h5F28207C;
    'h064B: mem_data <= 32'h207C2029;
    'h064C: mem_data <= 32'h5F5F5F7C;
    'h064D: mem_data <= 32'h0000000A;
    'h064E: mem_data <= 32'h7C5F7C20;
    'h064F: mem_data <= 32'h7C202020;
    'h0650: mem_data <= 32'h5F5C7C5F;
    'h0651: mem_data <= 32'h5F5C5F5F;
    'h0652: mem_data <= 32'h5F2F5F5F;
    'h0653: mem_data <= 32'h2F5F5F5F;
    'h0654: mem_data <= 32'h5F5F5C20;
    'h0655: mem_data <= 32'h5C202F5F;
    'h0656: mem_data <= 32'h5F5F5F5F;
    'h0657: mem_data <= 32'h00000A7C;
    'h0658: mem_data <= 32'h20495053;
    'h0659: mem_data <= 32'h74617453;
    'h065A: mem_data <= 32'h000A3A65;
    'h065B: mem_data <= 32'h414C2020;
    'h065C: mem_data <= 32'h434E4554;
    'h065D: mem_data <= 32'h00002059;
    'h065E: mem_data <= 32'h44442020;
    'h065F: mem_data <= 32'h00002052;
    'h0660: mem_data <= 32'h000A4E4F;
    'h0661: mem_data <= 32'h0A46464F;
    'h0662: mem_data <= 32'h00000000;
    'h0663: mem_data <= 32'h53512020;
    'h0664: mem_data <= 32'h00204950;
    'h0665: mem_data <= 32'h52432020;
    'h0666: mem_data <= 32'h0000204D;
    'h0667: mem_data <= 32'h656C6553;
    'h0668: mem_data <= 32'h61207463;
    'h0669: mem_data <= 32'h6361206E;
    'h066A: mem_data <= 32'h6E6F6974;
    'h066B: mem_data <= 32'h00000A3A;
    'h066C: mem_data <= 32'h5B202020;
    'h066D: mem_data <= 32'h52205D31;
    'h066E: mem_data <= 32'h20646165;
    'h066F: mem_data <= 32'h20495053;
    'h0670: mem_data <= 32'h73616C46;
    'h0671: mem_data <= 32'h44492068;
    'h0672: mem_data <= 32'h0000000A;
    'h0673: mem_data <= 32'h5B202020;
    'h0674: mem_data <= 32'h52205D32;
    'h0675: mem_data <= 32'h20646165;
    'h0676: mem_data <= 32'h20495053;
    'h0677: mem_data <= 32'h666E6F43;
    'h0678: mem_data <= 32'h52206769;
    'h0679: mem_data <= 32'h0A736765;
    'h067A: mem_data <= 32'h00000000;
    'h067B: mem_data <= 32'h5B202020;
    'h067C: mem_data <= 32'h53205D33;
    'h067D: mem_data <= 32'h63746977;
    'h067E: mem_data <= 32'h6F742068;
    'h067F: mem_data <= 32'h66656420;
    'h0680: mem_data <= 32'h746C7561;
    'h0681: mem_data <= 32'h646F6D20;
    'h0682: mem_data <= 32'h00000A65;
    'h0683: mem_data <= 32'h5B202020;
    'h0684: mem_data <= 32'h53205D34;
    'h0685: mem_data <= 32'h63746977;
    'h0686: mem_data <= 32'h6F742068;
    'h0687: mem_data <= 32'h61754420;
    'h0688: mem_data <= 32'h2F49206C;
    'h0689: mem_data <= 32'h6F6D204F;
    'h068A: mem_data <= 32'h000A6564;
    'h068B: mem_data <= 32'h5B202020;
    'h068C: mem_data <= 32'h53205D35;
    'h068D: mem_data <= 32'h63746977;
    'h068E: mem_data <= 32'h6F742068;
    'h068F: mem_data <= 32'h61755120;
    'h0690: mem_data <= 32'h2F492064;
    'h0691: mem_data <= 32'h6F6D204F;
    'h0692: mem_data <= 32'h000A6564;
    'h0693: mem_data <= 32'h5B202020;
    'h0694: mem_data <= 32'h53205D36;
    'h0695: mem_data <= 32'h63746977;
    'h0696: mem_data <= 32'h6F742068;
    'h0697: mem_data <= 32'h61755120;
    'h0698: mem_data <= 32'h44442064;
    'h0699: mem_data <= 32'h6F6D2052;
    'h069A: mem_data <= 32'h000A6564;
    'h069B: mem_data <= 32'h5B202020;
    'h069C: mem_data <= 32'h54205D37;
    'h069D: mem_data <= 32'h6C67676F;
    'h069E: mem_data <= 32'h6F632065;
    'h069F: mem_data <= 32'h6E69746E;
    'h06A0: mem_data <= 32'h73756F75;
    'h06A1: mem_data <= 32'h61657220;
    'h06A2: mem_data <= 32'h6F6D2064;
    'h06A3: mem_data <= 32'h000A6564;
    'h06A4: mem_data <= 32'h5B202020;
    'h06A5: mem_data <= 32'h52205D39;
    'h06A6: mem_data <= 32'h73206E75;
    'h06A7: mem_data <= 32'h6C706D69;
    'h06A8: mem_data <= 32'h69747369;
    'h06A9: mem_data <= 32'h65622063;
    'h06AA: mem_data <= 32'h6D68636E;
    'h06AB: mem_data <= 32'h0A6B7261;
    'h06AC: mem_data <= 32'h00000000;
    'h06AD: mem_data <= 32'h5B202020;
    'h06AE: mem_data <= 32'h42205D30;
    'h06AF: mem_data <= 32'h68636E65;
    'h06B0: mem_data <= 32'h6B72616D;
    'h06B1: mem_data <= 32'h6C6C6120;
    'h06B2: mem_data <= 32'h6E6F6320;
    'h06B3: mem_data <= 32'h73676966;
    'h06B4: mem_data <= 32'h0000000A;
    'h06B5: mem_data <= 32'h6D6D6F43;
    'h06B6: mem_data <= 32'h3E646E61;
    'h06B7: mem_data <= 32'h00000020;
    'h06B8: mem_data <= 32'h0010174C;
    'h06B9: mem_data <= 32'h001016F0;
    'h06BA: mem_data <= 32'h001016F8;
    'h06BB: mem_data <= 32'h00101700;
    'h06BC: mem_data <= 32'h00101708;
    'h06BD: mem_data <= 32'h00101710;
    'h06BE: mem_data <= 32'h00101718;
    'h06BF: mem_data <= 32'h00101720;
    'h06C0: mem_data <= 32'h00101754;
    'h06C1: mem_data <= 32'h0010173C;


    default:    mem_data <= 32'hDEADBEEF;

    endcase

// ============================================================================

reg o_ready;

always @(posedge clk or negedge rstn)
    if (!rstn)  o_ready <= 1'd0;
    else        o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

// Output connectins
assign ready    = o_ready;
assign rdata    = mem_data;
assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule
